LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

entity d8m_gpio is
	port (
		clk: in std_logic 
	);
end entity;
