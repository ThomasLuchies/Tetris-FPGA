-- sram.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sram is
	port (
		clk_clk             : in    std_logic                     := '0';             --          clk.clk
		hex7_export         : out   std_logic_vector(6 downto 0);                     --         hex7.export
		hex_0_export        : out   std_logic_vector(6 downto 0);                     --        hex_0.export
		hex_1_export        : out   std_logic_vector(6 downto 0);                     --        hex_1.export
		hex_2_export        : out   std_logic_vector(6 downto 0);                     --        hex_2.export
		hex_3_export        : out   std_logic_vector(6 downto 0);                     --        hex_3.export
		hex_4_export        : out   std_logic_vector(6 downto 0);                     --        hex_4.export
		hex_5_export        : out   std_logic_vector(6 downto 0);                     --        hex_5.export
		hex_6_export        : out   std_logic_vector(6 downto 0);                     --        hex_6.export
		move_left_export    : in    std_logic                     := '0';             --    move_left.export
		move_right_export   : in    std_logic                     := '0';             --   move_right.export
		reset_reset_n       : in    std_logic                     := '0';             --        reset.reset_n
		rotate_left_export  : in    std_logic                     := '0';             --  rotate_left.export
		rotate_right_export : in    std_logic                     := '0';             -- rotate_right.export
		row_0_export        : out   std_logic_vector(29 downto 0);                    --        row_0.export
		row_1_export        : out   std_logic_vector(29 downto 0);                    --        row_1.export
		row_10_export       : out   std_logic_vector(29 downto 0);                    --       row_10.export
		row_11_export       : out   std_logic_vector(29 downto 0);                    --       row_11.export
		row_12_export       : out   std_logic_vector(29 downto 0);                    --       row_12.export
		row_13_export       : out   std_logic_vector(29 downto 0);                    --       row_13.export
		row_14_export       : out   std_logic_vector(29 downto 0);                    --       row_14.export
		row_15_export       : out   std_logic_vector(29 downto 0);                    --       row_15.export
		row_16_export       : out   std_logic_vector(29 downto 0);                    --       row_16.export
		row_17_export       : out   std_logic_vector(29 downto 0);                    --       row_17.export
		row_18_export       : out   std_logic_vector(29 downto 0);                    --       row_18.export
		row_19_export       : out   std_logic_vector(29 downto 0);                    --       row_19.export
		row_2_export        : out   std_logic_vector(29 downto 0);                    --        row_2.export
		row_20_export       : out   std_logic_vector(29 downto 0);                    --       row_20.export
		row_21_export       : out   std_logic_vector(29 downto 0);                    --       row_21.export
		row_22_export       : out   std_logic_vector(29 downto 0);                    --       row_22.export
		row_23_export       : out   std_logic_vector(29 downto 0);                    --       row_23.export
		row_3_export        : out   std_logic_vector(29 downto 0);                    --        row_3.export
		row_4_export        : out   std_logic_vector(29 downto 0);                    --        row_4.export
		row_5_export        : out   std_logic_vector(29 downto 0);                    --        row_5.export
		row_6_export        : out   std_logic_vector(29 downto 0);                    --        row_6.export
		row_7_export        : out   std_logic_vector(29 downto 0);                    --        row_7.export
		row_8_export        : out   std_logic_vector(29 downto 0);                    --        row_8.export
		row_9_export        : out   std_logic_vector(29 downto 0);                    --        row_9.export
		sram_DQ             : inout std_logic_vector(15 downto 0) := (others => '0'); --         sram.DQ
		sram_ADDR           : out   std_logic_vector(19 downto 0);                    --             .ADDR
		sram_LB_N           : out   std_logic;                                        --             .LB_N
		sram_UB_N           : out   std_logic;                                        --             .UB_N
		sram_CE_N           : out   std_logic;                                        --             .CE_N
		sram_OE_N           : out   std_logic;                                        --             .OE_N
		sram_WE_N           : out   std_logic                                         --             .WE_N
	);
end entity sram;

architecture rtl of sram is
	component sram_HEX_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component sram_HEX_0;

	component sram_frame_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component sram_frame_timer;

	component sram_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component sram_jtag_uart_0;

	component sram_move_left is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component sram_move_left;

	component sram_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(25 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(21 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component sram_nios2_gen2_0;

	component sram_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component sram_onchip_memory2_0;

	component sram_row_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(29 downto 0)                     -- export
		);
	end component sram_row_0;

	component sram_sram_0 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component sram_sram_0;

	component sram_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address               : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address        : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			frame_timer_s1_address                         : out std_logic_vector(2 downto 0);                     -- address
			frame_timer_s1_write                           : out std_logic;                                        -- write
			frame_timer_s1_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			frame_timer_s1_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			frame_timer_s1_chipselect                      : out std_logic;                                        -- chipselect
			HEX_0_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			HEX_0_s1_write                                 : out std_logic;                                        -- write
			HEX_0_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_0_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_0_s1_chipselect                            : out std_logic;                                        -- chipselect
			HEX_1_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			HEX_1_s1_write                                 : out std_logic;                                        -- write
			HEX_1_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_1_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_1_s1_chipselect                            : out std_logic;                                        -- chipselect
			HEX_2_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			HEX_2_s1_write                                 : out std_logic;                                        -- write
			HEX_2_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_2_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_2_s1_chipselect                            : out std_logic;                                        -- chipselect
			HEX_3_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			HEX_3_s1_write                                 : out std_logic;                                        -- write
			HEX_3_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_3_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_3_s1_chipselect                            : out std_logic;                                        -- chipselect
			HEX_4_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			HEX_4_s1_write                                 : out std_logic;                                        -- write
			HEX_4_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_4_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_4_s1_chipselect                            : out std_logic;                                        -- chipselect
			HEX_5_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			HEX_5_s1_write                                 : out std_logic;                                        -- write
			HEX_5_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_5_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_5_s1_chipselect                            : out std_logic;                                        -- chipselect
			HEX_6_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			HEX_6_s1_write                                 : out std_logic;                                        -- write
			HEX_6_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_6_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_6_s1_chipselect                            : out std_logic;                                        -- chipselect
			HEX_7_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			HEX_7_s1_write                                 : out std_logic;                                        -- write
			HEX_7_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_7_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_7_s1_chipselect                            : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write            : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read             : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			move_left_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			move_left_s1_write                             : out std_logic;                                        -- write
			move_left_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			move_left_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			move_left_s1_chipselect                        : out std_logic;                                        -- chipselect
			move_right_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			move_right_s1_write                            : out std_logic;                                        -- write
			move_right_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			move_right_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			move_right_s1_chipselect                       : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                    : out std_logic_vector(16 downto 0);                    -- address
			onchip_memory2_0_s1_write                      : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                  : out std_logic_vector(15 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                 : out std_logic_vector(1 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                 : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                      : out std_logic;                                        -- clken
			rotate_left_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			rotate_left_s1_write                           : out std_logic;                                        -- write
			rotate_left_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rotate_left_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			rotate_left_s1_chipselect                      : out std_logic;                                        -- chipselect
			rotate_right_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			rotate_right_s1_write                          : out std_logic;                                        -- write
			rotate_right_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rotate_right_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			rotate_right_s1_chipselect                     : out std_logic;                                        -- chipselect
			row_0_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_0_s1_write                                 : out std_logic;                                        -- write
			row_0_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_0_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_0_s1_chipselect                            : out std_logic;                                        -- chipselect
			row_1_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_1_s1_write                                 : out std_logic;                                        -- write
			row_1_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_1_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_1_s1_chipselect                            : out std_logic;                                        -- chipselect
			row_10_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_10_s1_write                                : out std_logic;                                        -- write
			row_10_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_10_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_10_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_11_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_11_s1_write                                : out std_logic;                                        -- write
			row_11_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_11_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_11_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_12_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_12_s1_write                                : out std_logic;                                        -- write
			row_12_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_12_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_12_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_13_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_13_s1_write                                : out std_logic;                                        -- write
			row_13_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_13_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_13_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_14_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_14_s1_write                                : out std_logic;                                        -- write
			row_14_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_14_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_14_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_15_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_15_s1_write                                : out std_logic;                                        -- write
			row_15_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_15_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_15_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_16_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_16_s1_write                                : out std_logic;                                        -- write
			row_16_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_16_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_16_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_17_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_17_s1_write                                : out std_logic;                                        -- write
			row_17_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_17_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_17_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_18_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_18_s1_write                                : out std_logic;                                        -- write
			row_18_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_18_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_18_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_19_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_19_s1_write                                : out std_logic;                                        -- write
			row_19_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_19_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_19_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_2_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_2_s1_write                                 : out std_logic;                                        -- write
			row_2_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_2_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_2_s1_chipselect                            : out std_logic;                                        -- chipselect
			row_20_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_20_s1_write                                : out std_logic;                                        -- write
			row_20_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_20_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_20_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_21_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_21_s1_write                                : out std_logic;                                        -- write
			row_21_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_21_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_21_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_22_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_22_s1_write                                : out std_logic;                                        -- write
			row_22_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_22_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_22_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_23_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			row_23_s1_write                                : out std_logic;                                        -- write
			row_23_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_23_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			row_23_s1_chipselect                           : out std_logic;                                        -- chipselect
			row_3_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_3_s1_write                                 : out std_logic;                                        -- write
			row_3_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_3_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_3_s1_chipselect                            : out std_logic;                                        -- chipselect
			row_4_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_4_s1_write                                 : out std_logic;                                        -- write
			row_4_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_4_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_4_s1_chipselect                            : out std_logic;                                        -- chipselect
			row_5_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_5_s1_write                                 : out std_logic;                                        -- write
			row_5_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_5_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_5_s1_chipselect                            : out std_logic;                                        -- chipselect
			row_6_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_6_s1_write                                 : out std_logic;                                        -- write
			row_6_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_6_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_6_s1_chipselect                            : out std_logic;                                        -- chipselect
			row_7_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_7_s1_write                                 : out std_logic;                                        -- write
			row_7_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_7_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_7_s1_chipselect                            : out std_logic;                                        -- chipselect
			row_8_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_8_s1_write                                 : out std_logic;                                        -- write
			row_8_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_8_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_8_s1_chipselect                            : out std_logic;                                        -- chipselect
			row_9_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			row_9_s1_write                                 : out std_logic;                                        -- write
			row_9_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			row_9_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			row_9_s1_chipselect                            : out std_logic;                                        -- chipselect
			sram_0_avalon_sram_slave_address               : out std_logic_vector(19 downto 0);                    -- address
			sram_0_avalon_sram_slave_write                 : out std_logic;                                        -- write
			sram_0_avalon_sram_slave_read                  : out std_logic;                                        -- read
			sram_0_avalon_sram_slave_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sram_0_avalon_sram_slave_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			sram_0_avalon_sram_slave_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			sram_0_avalon_sram_slave_readdatavalid         : in  std_logic                     := 'X'              -- readdatavalid
		);
	end component sram_mm_interconnect_0;

	component sram_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component sram_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_gen2_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                            : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                : std_logic_vector(25 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                   : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                  : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                         : std_logic_vector(21 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                            : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sram_0_avalon_sram_slave_readdata             : std_logic_vector(15 downto 0); -- sram_0:readdata -> mm_interconnect_0:sram_0_avalon_sram_slave_readdata
	signal mm_interconnect_0_sram_0_avalon_sram_slave_address              : std_logic_vector(19 downto 0); -- mm_interconnect_0:sram_0_avalon_sram_slave_address -> sram_0:address
	signal mm_interconnect_0_sram_0_avalon_sram_slave_read                 : std_logic;                     -- mm_interconnect_0:sram_0_avalon_sram_slave_read -> sram_0:read
	signal mm_interconnect_0_sram_0_avalon_sram_slave_byteenable           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sram_0_avalon_sram_slave_byteenable -> sram_0:byteenable
	signal mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid        : std_logic;                     -- sram_0:readdatavalid -> mm_interconnect_0:sram_0_avalon_sram_slave_readdatavalid
	signal mm_interconnect_0_sram_0_avalon_sram_slave_write                : std_logic;                     -- mm_interconnect_0:sram_0_avalon_sram_slave_write -> sram_0:write
	signal mm_interconnect_0_sram_0_avalon_sram_slave_writedata            : std_logic_vector(15 downto 0); -- mm_interconnect_0:sram_0_avalon_sram_slave_writedata -> sram_0:writedata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                  : std_logic_vector(15 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                   : std_logic_vector(16 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_row_0_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_0_s1_chipselect -> row_0:chipselect
	signal mm_interconnect_0_row_0_s1_readdata                             : std_logic_vector(31 downto 0); -- row_0:readdata -> mm_interconnect_0:row_0_s1_readdata
	signal mm_interconnect_0_row_0_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_0_s1_address -> row_0:address
	signal mm_interconnect_0_row_0_s1_write                                : std_logic;                     -- mm_interconnect_0:row_0_s1_write -> mm_interconnect_0_row_0_s1_write:in
	signal mm_interconnect_0_row_0_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_0_s1_writedata -> row_0:writedata
	signal mm_interconnect_0_row_1_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_1_s1_chipselect -> row_1:chipselect
	signal mm_interconnect_0_row_1_s1_readdata                             : std_logic_vector(31 downto 0); -- row_1:readdata -> mm_interconnect_0:row_1_s1_readdata
	signal mm_interconnect_0_row_1_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_1_s1_address -> row_1:address
	signal mm_interconnect_0_row_1_s1_write                                : std_logic;                     -- mm_interconnect_0:row_1_s1_write -> mm_interconnect_0_row_1_s1_write:in
	signal mm_interconnect_0_row_1_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_1_s1_writedata -> row_1:writedata
	signal mm_interconnect_0_row_2_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_2_s1_chipselect -> row_2:chipselect
	signal mm_interconnect_0_row_2_s1_readdata                             : std_logic_vector(31 downto 0); -- row_2:readdata -> mm_interconnect_0:row_2_s1_readdata
	signal mm_interconnect_0_row_2_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_2_s1_address -> row_2:address
	signal mm_interconnect_0_row_2_s1_write                                : std_logic;                     -- mm_interconnect_0:row_2_s1_write -> mm_interconnect_0_row_2_s1_write:in
	signal mm_interconnect_0_row_2_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_2_s1_writedata -> row_2:writedata
	signal mm_interconnect_0_row_3_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_3_s1_chipselect -> row_3:chipselect
	signal mm_interconnect_0_row_3_s1_readdata                             : std_logic_vector(31 downto 0); -- row_3:readdata -> mm_interconnect_0:row_3_s1_readdata
	signal mm_interconnect_0_row_3_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_3_s1_address -> row_3:address
	signal mm_interconnect_0_row_3_s1_write                                : std_logic;                     -- mm_interconnect_0:row_3_s1_write -> mm_interconnect_0_row_3_s1_write:in
	signal mm_interconnect_0_row_3_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_3_s1_writedata -> row_3:writedata
	signal mm_interconnect_0_row_4_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_4_s1_chipselect -> row_4:chipselect
	signal mm_interconnect_0_row_4_s1_readdata                             : std_logic_vector(31 downto 0); -- row_4:readdata -> mm_interconnect_0:row_4_s1_readdata
	signal mm_interconnect_0_row_4_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_4_s1_address -> row_4:address
	signal mm_interconnect_0_row_4_s1_write                                : std_logic;                     -- mm_interconnect_0:row_4_s1_write -> mm_interconnect_0_row_4_s1_write:in
	signal mm_interconnect_0_row_4_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_4_s1_writedata -> row_4:writedata
	signal mm_interconnect_0_row_5_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_5_s1_chipselect -> row_5:chipselect
	signal mm_interconnect_0_row_5_s1_readdata                             : std_logic_vector(31 downto 0); -- row_5:readdata -> mm_interconnect_0:row_5_s1_readdata
	signal mm_interconnect_0_row_5_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_5_s1_address -> row_5:address
	signal mm_interconnect_0_row_5_s1_write                                : std_logic;                     -- mm_interconnect_0:row_5_s1_write -> mm_interconnect_0_row_5_s1_write:in
	signal mm_interconnect_0_row_5_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_5_s1_writedata -> row_5:writedata
	signal mm_interconnect_0_row_6_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_6_s1_chipselect -> row_6:chipselect
	signal mm_interconnect_0_row_6_s1_readdata                             : std_logic_vector(31 downto 0); -- row_6:readdata -> mm_interconnect_0:row_6_s1_readdata
	signal mm_interconnect_0_row_6_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_6_s1_address -> row_6:address
	signal mm_interconnect_0_row_6_s1_write                                : std_logic;                     -- mm_interconnect_0:row_6_s1_write -> mm_interconnect_0_row_6_s1_write:in
	signal mm_interconnect_0_row_6_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_6_s1_writedata -> row_6:writedata
	signal mm_interconnect_0_row_7_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_7_s1_chipselect -> row_7:chipselect
	signal mm_interconnect_0_row_7_s1_readdata                             : std_logic_vector(31 downto 0); -- row_7:readdata -> mm_interconnect_0:row_7_s1_readdata
	signal mm_interconnect_0_row_7_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_7_s1_address -> row_7:address
	signal mm_interconnect_0_row_7_s1_write                                : std_logic;                     -- mm_interconnect_0:row_7_s1_write -> mm_interconnect_0_row_7_s1_write:in
	signal mm_interconnect_0_row_7_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_7_s1_writedata -> row_7:writedata
	signal mm_interconnect_0_row_8_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_8_s1_chipselect -> row_8:chipselect
	signal mm_interconnect_0_row_8_s1_readdata                             : std_logic_vector(31 downto 0); -- row_8:readdata -> mm_interconnect_0:row_8_s1_readdata
	signal mm_interconnect_0_row_8_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_8_s1_address -> row_8:address
	signal mm_interconnect_0_row_8_s1_write                                : std_logic;                     -- mm_interconnect_0:row_8_s1_write -> mm_interconnect_0_row_8_s1_write:in
	signal mm_interconnect_0_row_8_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_8_s1_writedata -> row_8:writedata
	signal mm_interconnect_0_row_9_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:row_9_s1_chipselect -> row_9:chipselect
	signal mm_interconnect_0_row_9_s1_readdata                             : std_logic_vector(31 downto 0); -- row_9:readdata -> mm_interconnect_0:row_9_s1_readdata
	signal mm_interconnect_0_row_9_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_9_s1_address -> row_9:address
	signal mm_interconnect_0_row_9_s1_write                                : std_logic;                     -- mm_interconnect_0:row_9_s1_write -> mm_interconnect_0_row_9_s1_write:in
	signal mm_interconnect_0_row_9_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_9_s1_writedata -> row_9:writedata
	signal mm_interconnect_0_row_11_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_11_s1_chipselect -> row_11:chipselect
	signal mm_interconnect_0_row_11_s1_readdata                            : std_logic_vector(31 downto 0); -- row_11:readdata -> mm_interconnect_0:row_11_s1_readdata
	signal mm_interconnect_0_row_11_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_11_s1_address -> row_11:address
	signal mm_interconnect_0_row_11_s1_write                               : std_logic;                     -- mm_interconnect_0:row_11_s1_write -> mm_interconnect_0_row_11_s1_write:in
	signal mm_interconnect_0_row_11_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_11_s1_writedata -> row_11:writedata
	signal mm_interconnect_0_row_12_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_12_s1_chipselect -> row_12:chipselect
	signal mm_interconnect_0_row_12_s1_readdata                            : std_logic_vector(31 downto 0); -- row_12:readdata -> mm_interconnect_0:row_12_s1_readdata
	signal mm_interconnect_0_row_12_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_12_s1_address -> row_12:address
	signal mm_interconnect_0_row_12_s1_write                               : std_logic;                     -- mm_interconnect_0:row_12_s1_write -> mm_interconnect_0_row_12_s1_write:in
	signal mm_interconnect_0_row_12_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_12_s1_writedata -> row_12:writedata
	signal mm_interconnect_0_row_13_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_13_s1_chipselect -> row_13:chipselect
	signal mm_interconnect_0_row_13_s1_readdata                            : std_logic_vector(31 downto 0); -- row_13:readdata -> mm_interconnect_0:row_13_s1_readdata
	signal mm_interconnect_0_row_13_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_13_s1_address -> row_13:address
	signal mm_interconnect_0_row_13_s1_write                               : std_logic;                     -- mm_interconnect_0:row_13_s1_write -> mm_interconnect_0_row_13_s1_write:in
	signal mm_interconnect_0_row_13_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_13_s1_writedata -> row_13:writedata
	signal mm_interconnect_0_row_14_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_14_s1_chipselect -> row_14:chipselect
	signal mm_interconnect_0_row_14_s1_readdata                            : std_logic_vector(31 downto 0); -- row_14:readdata -> mm_interconnect_0:row_14_s1_readdata
	signal mm_interconnect_0_row_14_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_14_s1_address -> row_14:address
	signal mm_interconnect_0_row_14_s1_write                               : std_logic;                     -- mm_interconnect_0:row_14_s1_write -> mm_interconnect_0_row_14_s1_write:in
	signal mm_interconnect_0_row_14_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_14_s1_writedata -> row_14:writedata
	signal mm_interconnect_0_row_15_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_15_s1_chipselect -> row_15:chipselect
	signal mm_interconnect_0_row_15_s1_readdata                            : std_logic_vector(31 downto 0); -- row_15:readdata -> mm_interconnect_0:row_15_s1_readdata
	signal mm_interconnect_0_row_15_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_15_s1_address -> row_15:address
	signal mm_interconnect_0_row_15_s1_write                               : std_logic;                     -- mm_interconnect_0:row_15_s1_write -> mm_interconnect_0_row_15_s1_write:in
	signal mm_interconnect_0_row_15_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_15_s1_writedata -> row_15:writedata
	signal mm_interconnect_0_row_16_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_16_s1_chipselect -> row_16:chipselect
	signal mm_interconnect_0_row_16_s1_readdata                            : std_logic_vector(31 downto 0); -- row_16:readdata -> mm_interconnect_0:row_16_s1_readdata
	signal mm_interconnect_0_row_16_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_16_s1_address -> row_16:address
	signal mm_interconnect_0_row_16_s1_write                               : std_logic;                     -- mm_interconnect_0:row_16_s1_write -> mm_interconnect_0_row_16_s1_write:in
	signal mm_interconnect_0_row_16_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_16_s1_writedata -> row_16:writedata
	signal mm_interconnect_0_row_17_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_17_s1_chipselect -> row_17:chipselect
	signal mm_interconnect_0_row_17_s1_readdata                            : std_logic_vector(31 downto 0); -- row_17:readdata -> mm_interconnect_0:row_17_s1_readdata
	signal mm_interconnect_0_row_17_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_17_s1_address -> row_17:address
	signal mm_interconnect_0_row_17_s1_write                               : std_logic;                     -- mm_interconnect_0:row_17_s1_write -> mm_interconnect_0_row_17_s1_write:in
	signal mm_interconnect_0_row_17_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_17_s1_writedata -> row_17:writedata
	signal mm_interconnect_0_row_18_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_18_s1_chipselect -> row_18:chipselect
	signal mm_interconnect_0_row_18_s1_readdata                            : std_logic_vector(31 downto 0); -- row_18:readdata -> mm_interconnect_0:row_18_s1_readdata
	signal mm_interconnect_0_row_18_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_18_s1_address -> row_18:address
	signal mm_interconnect_0_row_18_s1_write                               : std_logic;                     -- mm_interconnect_0:row_18_s1_write -> mm_interconnect_0_row_18_s1_write:in
	signal mm_interconnect_0_row_18_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_18_s1_writedata -> row_18:writedata
	signal mm_interconnect_0_row_19_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_19_s1_chipselect -> row_19:chipselect
	signal mm_interconnect_0_row_19_s1_readdata                            : std_logic_vector(31 downto 0); -- row_19:readdata -> mm_interconnect_0:row_19_s1_readdata
	signal mm_interconnect_0_row_19_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_19_s1_address -> row_19:address
	signal mm_interconnect_0_row_19_s1_write                               : std_logic;                     -- mm_interconnect_0:row_19_s1_write -> mm_interconnect_0_row_19_s1_write:in
	signal mm_interconnect_0_row_19_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_19_s1_writedata -> row_19:writedata
	signal mm_interconnect_0_row_20_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_20_s1_chipselect -> row_20:chipselect
	signal mm_interconnect_0_row_20_s1_readdata                            : std_logic_vector(31 downto 0); -- row_20:readdata -> mm_interconnect_0:row_20_s1_readdata
	signal mm_interconnect_0_row_20_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_20_s1_address -> row_20:address
	signal mm_interconnect_0_row_20_s1_write                               : std_logic;                     -- mm_interconnect_0:row_20_s1_write -> mm_interconnect_0_row_20_s1_write:in
	signal mm_interconnect_0_row_20_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_20_s1_writedata -> row_20:writedata
	signal mm_interconnect_0_row_21_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_21_s1_chipselect -> row_21:chipselect
	signal mm_interconnect_0_row_21_s1_readdata                            : std_logic_vector(31 downto 0); -- row_21:readdata -> mm_interconnect_0:row_21_s1_readdata
	signal mm_interconnect_0_row_21_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_21_s1_address -> row_21:address
	signal mm_interconnect_0_row_21_s1_write                               : std_logic;                     -- mm_interconnect_0:row_21_s1_write -> mm_interconnect_0_row_21_s1_write:in
	signal mm_interconnect_0_row_21_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_21_s1_writedata -> row_21:writedata
	signal mm_interconnect_0_row_22_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_22_s1_chipselect -> row_22:chipselect
	signal mm_interconnect_0_row_22_s1_readdata                            : std_logic_vector(31 downto 0); -- row_22:readdata -> mm_interconnect_0:row_22_s1_readdata
	signal mm_interconnect_0_row_22_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_22_s1_address -> row_22:address
	signal mm_interconnect_0_row_22_s1_write                               : std_logic;                     -- mm_interconnect_0:row_22_s1_write -> mm_interconnect_0_row_22_s1_write:in
	signal mm_interconnect_0_row_22_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_22_s1_writedata -> row_22:writedata
	signal mm_interconnect_0_row_23_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_23_s1_chipselect -> row_23:chipselect
	signal mm_interconnect_0_row_23_s1_readdata                            : std_logic_vector(31 downto 0); -- row_23:readdata -> mm_interconnect_0:row_23_s1_readdata
	signal mm_interconnect_0_row_23_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_23_s1_address -> row_23:address
	signal mm_interconnect_0_row_23_s1_write                               : std_logic;                     -- mm_interconnect_0:row_23_s1_write -> mm_interconnect_0_row_23_s1_write:in
	signal mm_interconnect_0_row_23_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_23_s1_writedata -> row_23:writedata
	signal mm_interconnect_0_row_10_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:row_10_s1_chipselect -> row_10:chipselect
	signal mm_interconnect_0_row_10_s1_readdata                            : std_logic_vector(31 downto 0); -- row_10:readdata -> mm_interconnect_0:row_10_s1_readdata
	signal mm_interconnect_0_row_10_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:row_10_s1_address -> row_10:address
	signal mm_interconnect_0_row_10_s1_write                               : std_logic;                     -- mm_interconnect_0:row_10_s1_write -> mm_interconnect_0_row_10_s1_write:in
	signal mm_interconnect_0_row_10_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:row_10_s1_writedata -> row_10:writedata
	signal mm_interconnect_0_move_left_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:move_left_s1_chipselect -> move_left:chipselect
	signal mm_interconnect_0_move_left_s1_readdata                         : std_logic_vector(31 downto 0); -- move_left:readdata -> mm_interconnect_0:move_left_s1_readdata
	signal mm_interconnect_0_move_left_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:move_left_s1_address -> move_left:address
	signal mm_interconnect_0_move_left_s1_write                            : std_logic;                     -- mm_interconnect_0:move_left_s1_write -> mm_interconnect_0_move_left_s1_write:in
	signal mm_interconnect_0_move_left_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:move_left_s1_writedata -> move_left:writedata
	signal mm_interconnect_0_move_right_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:move_right_s1_chipselect -> move_right:chipselect
	signal mm_interconnect_0_move_right_s1_readdata                        : std_logic_vector(31 downto 0); -- move_right:readdata -> mm_interconnect_0:move_right_s1_readdata
	signal mm_interconnect_0_move_right_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:move_right_s1_address -> move_right:address
	signal mm_interconnect_0_move_right_s1_write                           : std_logic;                     -- mm_interconnect_0:move_right_s1_write -> mm_interconnect_0_move_right_s1_write:in
	signal mm_interconnect_0_move_right_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:move_right_s1_writedata -> move_right:writedata
	signal mm_interconnect_0_rotate_left_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:rotate_left_s1_chipselect -> rotate_left:chipselect
	signal mm_interconnect_0_rotate_left_s1_readdata                       : std_logic_vector(31 downto 0); -- rotate_left:readdata -> mm_interconnect_0:rotate_left_s1_readdata
	signal mm_interconnect_0_rotate_left_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:rotate_left_s1_address -> rotate_left:address
	signal mm_interconnect_0_rotate_left_s1_write                          : std_logic;                     -- mm_interconnect_0:rotate_left_s1_write -> mm_interconnect_0_rotate_left_s1_write:in
	signal mm_interconnect_0_rotate_left_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:rotate_left_s1_writedata -> rotate_left:writedata
	signal mm_interconnect_0_rotate_right_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:rotate_right_s1_chipselect -> rotate_right:chipselect
	signal mm_interconnect_0_rotate_right_s1_readdata                      : std_logic_vector(31 downto 0); -- rotate_right:readdata -> mm_interconnect_0:rotate_right_s1_readdata
	signal mm_interconnect_0_rotate_right_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:rotate_right_s1_address -> rotate_right:address
	signal mm_interconnect_0_rotate_right_s1_write                         : std_logic;                     -- mm_interconnect_0:rotate_right_s1_write -> mm_interconnect_0_rotate_right_s1_write:in
	signal mm_interconnect_0_rotate_right_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:rotate_right_s1_writedata -> rotate_right:writedata
	signal mm_interconnect_0_frame_timer_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:frame_timer_s1_chipselect -> frame_timer:chipselect
	signal mm_interconnect_0_frame_timer_s1_readdata                       : std_logic_vector(15 downto 0); -- frame_timer:readdata -> mm_interconnect_0:frame_timer_s1_readdata
	signal mm_interconnect_0_frame_timer_s1_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:frame_timer_s1_address -> frame_timer:address
	signal mm_interconnect_0_frame_timer_s1_write                          : std_logic;                     -- mm_interconnect_0:frame_timer_s1_write -> mm_interconnect_0_frame_timer_s1_write:in
	signal mm_interconnect_0_frame_timer_s1_writedata                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:frame_timer_s1_writedata -> frame_timer:writedata
	signal mm_interconnect_0_hex_0_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:HEX_0_s1_chipselect -> HEX_0:chipselect
	signal mm_interconnect_0_hex_0_s1_readdata                             : std_logic_vector(31 downto 0); -- HEX_0:readdata -> mm_interconnect_0:HEX_0_s1_readdata
	signal mm_interconnect_0_hex_0_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_0_s1_address -> HEX_0:address
	signal mm_interconnect_0_hex_0_s1_write                                : std_logic;                     -- mm_interconnect_0:HEX_0_s1_write -> mm_interconnect_0_hex_0_s1_write:in
	signal mm_interconnect_0_hex_0_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_0_s1_writedata -> HEX_0:writedata
	signal mm_interconnect_0_hex_1_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:HEX_1_s1_chipselect -> HEX_1:chipselect
	signal mm_interconnect_0_hex_1_s1_readdata                             : std_logic_vector(31 downto 0); -- HEX_1:readdata -> mm_interconnect_0:HEX_1_s1_readdata
	signal mm_interconnect_0_hex_1_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_1_s1_address -> HEX_1:address
	signal mm_interconnect_0_hex_1_s1_write                                : std_logic;                     -- mm_interconnect_0:HEX_1_s1_write -> mm_interconnect_0_hex_1_s1_write:in
	signal mm_interconnect_0_hex_1_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_1_s1_writedata -> HEX_1:writedata
	signal mm_interconnect_0_hex_2_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:HEX_2_s1_chipselect -> HEX_2:chipselect
	signal mm_interconnect_0_hex_2_s1_readdata                             : std_logic_vector(31 downto 0); -- HEX_2:readdata -> mm_interconnect_0:HEX_2_s1_readdata
	signal mm_interconnect_0_hex_2_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_2_s1_address -> HEX_2:address
	signal mm_interconnect_0_hex_2_s1_write                                : std_logic;                     -- mm_interconnect_0:HEX_2_s1_write -> mm_interconnect_0_hex_2_s1_write:in
	signal mm_interconnect_0_hex_2_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_2_s1_writedata -> HEX_2:writedata
	signal mm_interconnect_0_hex_3_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:HEX_3_s1_chipselect -> HEX_3:chipselect
	signal mm_interconnect_0_hex_3_s1_readdata                             : std_logic_vector(31 downto 0); -- HEX_3:readdata -> mm_interconnect_0:HEX_3_s1_readdata
	signal mm_interconnect_0_hex_3_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_3_s1_address -> HEX_3:address
	signal mm_interconnect_0_hex_3_s1_write                                : std_logic;                     -- mm_interconnect_0:HEX_3_s1_write -> mm_interconnect_0_hex_3_s1_write:in
	signal mm_interconnect_0_hex_3_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_3_s1_writedata -> HEX_3:writedata
	signal mm_interconnect_0_hex_4_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:HEX_4_s1_chipselect -> HEX_4:chipselect
	signal mm_interconnect_0_hex_4_s1_readdata                             : std_logic_vector(31 downto 0); -- HEX_4:readdata -> mm_interconnect_0:HEX_4_s1_readdata
	signal mm_interconnect_0_hex_4_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_4_s1_address -> HEX_4:address
	signal mm_interconnect_0_hex_4_s1_write                                : std_logic;                     -- mm_interconnect_0:HEX_4_s1_write -> mm_interconnect_0_hex_4_s1_write:in
	signal mm_interconnect_0_hex_4_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_4_s1_writedata -> HEX_4:writedata
	signal mm_interconnect_0_hex_5_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:HEX_5_s1_chipselect -> HEX_5:chipselect
	signal mm_interconnect_0_hex_5_s1_readdata                             : std_logic_vector(31 downto 0); -- HEX_5:readdata -> mm_interconnect_0:HEX_5_s1_readdata
	signal mm_interconnect_0_hex_5_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_5_s1_address -> HEX_5:address
	signal mm_interconnect_0_hex_5_s1_write                                : std_logic;                     -- mm_interconnect_0:HEX_5_s1_write -> mm_interconnect_0_hex_5_s1_write:in
	signal mm_interconnect_0_hex_5_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_5_s1_writedata -> HEX_5:writedata
	signal mm_interconnect_0_hex_6_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:HEX_6_s1_chipselect -> HEX_6:chipselect
	signal mm_interconnect_0_hex_6_s1_readdata                             : std_logic_vector(31 downto 0); -- HEX_6:readdata -> mm_interconnect_0:HEX_6_s1_readdata
	signal mm_interconnect_0_hex_6_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_6_s1_address -> HEX_6:address
	signal mm_interconnect_0_hex_6_s1_write                                : std_logic;                     -- mm_interconnect_0:HEX_6_s1_write -> mm_interconnect_0_hex_6_s1_write:in
	signal mm_interconnect_0_hex_6_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_6_s1_writedata -> HEX_6:writedata
	signal mm_interconnect_0_hex_7_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:HEX_7_s1_chipselect -> HEX_7:chipselect
	signal mm_interconnect_0_hex_7_s1_readdata                             : std_logic_vector(31 downto 0); -- HEX_7:readdata -> mm_interconnect_0:HEX_7_s1_readdata
	signal mm_interconnect_0_hex_7_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_7_s1_address -> HEX_7:address
	signal mm_interconnect_0_hex_7_s1_write                                : std_logic;                     -- mm_interconnect_0:HEX_7_s1_write -> mm_interconnect_0_hex_7_s1_write:in
	signal mm_interconnect_0_hex_7_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_7_s1_writedata -> HEX_7:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- move_left:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- move_right:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- rotate_left:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                        : std_logic;                     -- rotate_right:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                        : std_logic;                     -- frame_timer:irq -> irq_mapper:receiver5_irq
	signal nios2_gen2_0_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, sram_0:reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                          : std_logic;                     -- nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_row_0_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_0_s1_write:inv -> row_0:write_n
	signal mm_interconnect_0_row_1_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_1_s1_write:inv -> row_1:write_n
	signal mm_interconnect_0_row_2_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_2_s1_write:inv -> row_2:write_n
	signal mm_interconnect_0_row_3_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_3_s1_write:inv -> row_3:write_n
	signal mm_interconnect_0_row_4_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_4_s1_write:inv -> row_4:write_n
	signal mm_interconnect_0_row_5_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_5_s1_write:inv -> row_5:write_n
	signal mm_interconnect_0_row_6_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_6_s1_write:inv -> row_6:write_n
	signal mm_interconnect_0_row_7_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_7_s1_write:inv -> row_7:write_n
	signal mm_interconnect_0_row_8_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_8_s1_write:inv -> row_8:write_n
	signal mm_interconnect_0_row_9_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_row_9_s1_write:inv -> row_9:write_n
	signal mm_interconnect_0_row_11_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_11_s1_write:inv -> row_11:write_n
	signal mm_interconnect_0_row_12_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_12_s1_write:inv -> row_12:write_n
	signal mm_interconnect_0_row_13_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_13_s1_write:inv -> row_13:write_n
	signal mm_interconnect_0_row_14_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_14_s1_write:inv -> row_14:write_n
	signal mm_interconnect_0_row_15_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_15_s1_write:inv -> row_15:write_n
	signal mm_interconnect_0_row_16_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_16_s1_write:inv -> row_16:write_n
	signal mm_interconnect_0_row_17_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_17_s1_write:inv -> row_17:write_n
	signal mm_interconnect_0_row_18_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_18_s1_write:inv -> row_18:write_n
	signal mm_interconnect_0_row_19_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_19_s1_write:inv -> row_19:write_n
	signal mm_interconnect_0_row_20_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_20_s1_write:inv -> row_20:write_n
	signal mm_interconnect_0_row_21_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_21_s1_write:inv -> row_21:write_n
	signal mm_interconnect_0_row_22_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_22_s1_write:inv -> row_22:write_n
	signal mm_interconnect_0_row_23_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_23_s1_write:inv -> row_23:write_n
	signal mm_interconnect_0_row_10_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_row_10_s1_write:inv -> row_10:write_n
	signal mm_interconnect_0_move_left_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_move_left_s1_write:inv -> move_left:write_n
	signal mm_interconnect_0_move_right_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_move_right_s1_write:inv -> move_right:write_n
	signal mm_interconnect_0_rotate_left_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_rotate_left_s1_write:inv -> rotate_left:write_n
	signal mm_interconnect_0_rotate_right_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_rotate_right_s1_write:inv -> rotate_right:write_n
	signal mm_interconnect_0_frame_timer_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_frame_timer_s1_write:inv -> frame_timer:write_n
	signal mm_interconnect_0_hex_0_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hex_0_s1_write:inv -> HEX_0:write_n
	signal mm_interconnect_0_hex_1_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hex_1_s1_write:inv -> HEX_1:write_n
	signal mm_interconnect_0_hex_2_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hex_2_s1_write:inv -> HEX_2:write_n
	signal mm_interconnect_0_hex_3_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hex_3_s1_write:inv -> HEX_3:write_n
	signal mm_interconnect_0_hex_4_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hex_4_s1_write:inv -> HEX_4:write_n
	signal mm_interconnect_0_hex_5_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hex_5_s1_write:inv -> HEX_5:write_n
	signal mm_interconnect_0_hex_6_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hex_6_s1_write:inv -> HEX_6:write_n
	signal mm_interconnect_0_hex_7_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hex_7_s1_write:inv -> HEX_7:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [HEX_0:reset_n, HEX_1:reset_n, HEX_2:reset_n, HEX_3:reset_n, HEX_4:reset_n, HEX_5:reset_n, HEX_6:reset_n, HEX_7:reset_n, frame_timer:reset_n, jtag_uart_0:rst_n, move_left:reset_n, move_right:reset_n, nios2_gen2_0:reset_n, rotate_left:reset_n, rotate_right:reset_n, row_0:reset_n, row_10:reset_n, row_11:reset_n, row_12:reset_n, row_13:reset_n, row_14:reset_n, row_15:reset_n, row_16:reset_n, row_17:reset_n, row_18:reset_n, row_19:reset_n, row_1:reset_n, row_20:reset_n, row_21:reset_n, row_22:reset_n, row_23:reset_n, row_2:reset_n, row_3:reset_n, row_4:reset_n, row_5:reset_n, row_6:reset_n, row_7:reset_n, row_8:reset_n, row_9:reset_n]

begin

	hex_0 : component sram_HEX_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_0_s1_readdata,        --                    .readdata
			out_port   => hex_0_export                                -- external_connection.export
		);

	hex_1 : component sram_HEX_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_1_s1_readdata,        --                    .readdata
			out_port   => hex_1_export                                -- external_connection.export
		);

	hex_2 : component sram_HEX_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_2_s1_readdata,        --                    .readdata
			out_port   => hex_2_export                                -- external_connection.export
		);

	hex_3 : component sram_HEX_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_3_s1_readdata,        --                    .readdata
			out_port   => hex_3_export                                -- external_connection.export
		);

	hex_4 : component sram_HEX_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_4_s1_readdata,        --                    .readdata
			out_port   => hex_4_export                                -- external_connection.export
		);

	hex_5 : component sram_HEX_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_5_s1_readdata,        --                    .readdata
			out_port   => hex_5_export                                -- external_connection.export
		);

	hex_6 : component sram_HEX_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_6_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_6_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_6_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_6_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_6_s1_readdata,        --                    .readdata
			out_port   => hex_6_export                                -- external_connection.export
		);

	hex_7 : component sram_HEX_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_7_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_7_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_7_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_7_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_7_s1_readdata,        --                    .readdata
			out_port   => hex7_export                                 -- external_connection.export
		);

	frame_timer : component sram_frame_timer
		port map (
			clk        => clk_clk,                                          --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         -- reset.reset_n
			address    => mm_interconnect_0_frame_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_frame_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_frame_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_frame_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_frame_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver5_irq                          --   irq.irq
		);

	jtag_uart_0 : component sram_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	move_left : component sram_move_left
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_move_left_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_move_left_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_move_left_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_move_left_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_move_left_s1_readdata,        --                    .readdata
			in_port    => move_left_export,                               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                        --                 irq.irq
		);

	move_right : component sram_move_left
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_move_right_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_move_right_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_move_right_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_move_right_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_move_right_s1_readdata,        --                    .readdata
			in_port    => move_right_export,                               -- external_connection.export
			irq        => irq_mapper_receiver2_irq                         --                 irq.irq
		);

	nios2_gen2_0 : component sram_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component sram_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	rotate_left : component sram_move_left
		port map (
			clk        => clk_clk,                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_rotate_left_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_rotate_left_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_rotate_left_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_rotate_left_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_rotate_left_s1_readdata,        --                    .readdata
			in_port    => rotate_left_export,                               -- external_connection.export
			irq        => irq_mapper_receiver3_irq                          --                 irq.irq
		);

	rotate_right : component sram_move_left
		port map (
			clk        => clk_clk,                                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_rotate_right_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_rotate_right_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_rotate_right_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_rotate_right_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_rotate_right_s1_readdata,        --                    .readdata
			in_port    => rotate_right_export,                               -- external_connection.export
			irq        => irq_mapper_receiver4_irq                           --                 irq.irq
		);

	row_0 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_0_s1_readdata,        --                    .readdata
			out_port   => row_0_export                                -- external_connection.export
		);

	row_1 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_1_s1_readdata,        --                    .readdata
			out_port   => row_1_export                                -- external_connection.export
		);

	row_10 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_10_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_10_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_10_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_10_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_10_s1_readdata,        --                    .readdata
			out_port   => row_10_export                                -- external_connection.export
		);

	row_11 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_11_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_11_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_11_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_11_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_11_s1_readdata,        --                    .readdata
			out_port   => row_11_export                                -- external_connection.export
		);

	row_12 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_12_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_12_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_12_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_12_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_12_s1_readdata,        --                    .readdata
			out_port   => row_12_export                                -- external_connection.export
		);

	row_13 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_13_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_13_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_13_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_13_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_13_s1_readdata,        --                    .readdata
			out_port   => row_13_export                                -- external_connection.export
		);

	row_14 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_14_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_14_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_14_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_14_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_14_s1_readdata,        --                    .readdata
			out_port   => row_14_export                                -- external_connection.export
		);

	row_15 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_15_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_15_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_15_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_15_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_15_s1_readdata,        --                    .readdata
			out_port   => row_15_export                                -- external_connection.export
		);

	row_16 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_16_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_16_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_16_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_16_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_16_s1_readdata,        --                    .readdata
			out_port   => row_16_export                                -- external_connection.export
		);

	row_17 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_17_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_17_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_17_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_17_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_17_s1_readdata,        --                    .readdata
			out_port   => row_17_export                                -- external_connection.export
		);

	row_18 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_18_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_18_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_18_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_18_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_18_s1_readdata,        --                    .readdata
			out_port   => row_18_export                                -- external_connection.export
		);

	row_19 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_19_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_19_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_19_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_19_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_19_s1_readdata,        --                    .readdata
			out_port   => row_19_export                                -- external_connection.export
		);

	row_2 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_2_s1_readdata,        --                    .readdata
			out_port   => row_2_export                                -- external_connection.export
		);

	row_20 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_20_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_20_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_20_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_20_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_20_s1_readdata,        --                    .readdata
			out_port   => row_20_export                                -- external_connection.export
		);

	row_21 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_21_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_21_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_21_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_21_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_21_s1_readdata,        --                    .readdata
			out_port   => row_21_export                                -- external_connection.export
		);

	row_22 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_22_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_22_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_22_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_22_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_22_s1_readdata,        --                    .readdata
			out_port   => row_22_export                                -- external_connection.export
		);

	row_23 : component sram_row_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_row_23_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_23_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_23_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_23_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_23_s1_readdata,        --                    .readdata
			out_port   => row_23_export                                -- external_connection.export
		);

	row_3 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_3_s1_readdata,        --                    .readdata
			out_port   => row_3_export                                -- external_connection.export
		);

	row_4 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_4_s1_readdata,        --                    .readdata
			out_port   => row_4_export                                -- external_connection.export
		);

	row_5 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_5_s1_readdata,        --                    .readdata
			out_port   => row_5_export                                -- external_connection.export
		);

	row_6 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_6_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_6_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_6_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_6_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_6_s1_readdata,        --                    .readdata
			out_port   => row_6_export                                -- external_connection.export
		);

	row_7 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_7_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_7_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_7_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_7_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_7_s1_readdata,        --                    .readdata
			out_port   => row_7_export                                -- external_connection.export
		);

	row_8 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_8_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_8_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_8_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_8_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_8_s1_readdata,        --                    .readdata
			out_port   => row_8_export                                -- external_connection.export
		);

	row_9 : component sram_row_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_row_9_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_row_9_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_row_9_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_row_9_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_row_9_s1_readdata,        --                    .readdata
			out_port   => row_9_export                                -- external_connection.export
		);

	sram_0 : component sram_sram_0
		port map (
			clk           => clk_clk,                                                  --                clk.clk
			reset         => rst_controller_reset_out_reset,                           --              reset.reset
			SRAM_DQ       => sram_DQ,                                                  -- external_interface.export
			SRAM_ADDR     => sram_ADDR,                                                --                   .export
			SRAM_LB_N     => sram_LB_N,                                                --                   .export
			SRAM_UB_N     => sram_UB_N,                                                --                   .export
			SRAM_CE_N     => sram_CE_N,                                                --                   .export
			SRAM_OE_N     => sram_OE_N,                                                --                   .export
			SRAM_WE_N     => sram_WE_N,                                                --                   .export
			address       => mm_interconnect_0_sram_0_avalon_sram_slave_address,       --  avalon_sram_slave.address
			byteenable    => mm_interconnect_0_sram_0_avalon_sram_slave_byteenable,    --                   .byteenable
			read          => mm_interconnect_0_sram_0_avalon_sram_slave_read,          --                   .read
			write         => mm_interconnect_0_sram_0_avalon_sram_slave_write,         --                   .write
			writedata     => mm_interconnect_0_sram_0_avalon_sram_slave_writedata,     --                   .writedata
			readdata      => mm_interconnect_0_sram_0_avalon_sram_slave_readdata,      --                   .readdata
			readdatavalid => mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid  --                   .readdatavalid
		);

	mm_interconnect_0 : component sram_mm_interconnect_0
		port map (
			clk_0_clk_clk                                  => clk_clk,                                                     --                                clk_0_clk.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address               => nios2_gen2_0_data_master_address,                            --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest           => nios2_gen2_0_data_master_waitrequest,                        --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable            => nios2_gen2_0_data_master_byteenable,                         --                                         .byteenable
			nios2_gen2_0_data_master_read                  => nios2_gen2_0_data_master_read,                               --                                         .read
			nios2_gen2_0_data_master_readdata              => nios2_gen2_0_data_master_readdata,                           --                                         .readdata
			nios2_gen2_0_data_master_write                 => nios2_gen2_0_data_master_write,                              --                                         .write
			nios2_gen2_0_data_master_writedata             => nios2_gen2_0_data_master_writedata,                          --                                         .writedata
			nios2_gen2_0_data_master_debugaccess           => nios2_gen2_0_data_master_debugaccess,                        --                                         .debugaccess
			nios2_gen2_0_instruction_master_address        => nios2_gen2_0_instruction_master_address,                     --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest    => nios2_gen2_0_instruction_master_waitrequest,                 --                                         .waitrequest
			nios2_gen2_0_instruction_master_read           => nios2_gen2_0_instruction_master_read,                        --                                         .read
			nios2_gen2_0_instruction_master_readdata       => nios2_gen2_0_instruction_master_readdata,                    --                                         .readdata
			frame_timer_s1_address                         => mm_interconnect_0_frame_timer_s1_address,                    --                           frame_timer_s1.address
			frame_timer_s1_write                           => mm_interconnect_0_frame_timer_s1_write,                      --                                         .write
			frame_timer_s1_readdata                        => mm_interconnect_0_frame_timer_s1_readdata,                   --                                         .readdata
			frame_timer_s1_writedata                       => mm_interconnect_0_frame_timer_s1_writedata,                  --                                         .writedata
			frame_timer_s1_chipselect                      => mm_interconnect_0_frame_timer_s1_chipselect,                 --                                         .chipselect
			HEX_0_s1_address                               => mm_interconnect_0_hex_0_s1_address,                          --                                 HEX_0_s1.address
			HEX_0_s1_write                                 => mm_interconnect_0_hex_0_s1_write,                            --                                         .write
			HEX_0_s1_readdata                              => mm_interconnect_0_hex_0_s1_readdata,                         --                                         .readdata
			HEX_0_s1_writedata                             => mm_interconnect_0_hex_0_s1_writedata,                        --                                         .writedata
			HEX_0_s1_chipselect                            => mm_interconnect_0_hex_0_s1_chipselect,                       --                                         .chipselect
			HEX_1_s1_address                               => mm_interconnect_0_hex_1_s1_address,                          --                                 HEX_1_s1.address
			HEX_1_s1_write                                 => mm_interconnect_0_hex_1_s1_write,                            --                                         .write
			HEX_1_s1_readdata                              => mm_interconnect_0_hex_1_s1_readdata,                         --                                         .readdata
			HEX_1_s1_writedata                             => mm_interconnect_0_hex_1_s1_writedata,                        --                                         .writedata
			HEX_1_s1_chipselect                            => mm_interconnect_0_hex_1_s1_chipselect,                       --                                         .chipselect
			HEX_2_s1_address                               => mm_interconnect_0_hex_2_s1_address,                          --                                 HEX_2_s1.address
			HEX_2_s1_write                                 => mm_interconnect_0_hex_2_s1_write,                            --                                         .write
			HEX_2_s1_readdata                              => mm_interconnect_0_hex_2_s1_readdata,                         --                                         .readdata
			HEX_2_s1_writedata                             => mm_interconnect_0_hex_2_s1_writedata,                        --                                         .writedata
			HEX_2_s1_chipselect                            => mm_interconnect_0_hex_2_s1_chipselect,                       --                                         .chipselect
			HEX_3_s1_address                               => mm_interconnect_0_hex_3_s1_address,                          --                                 HEX_3_s1.address
			HEX_3_s1_write                                 => mm_interconnect_0_hex_3_s1_write,                            --                                         .write
			HEX_3_s1_readdata                              => mm_interconnect_0_hex_3_s1_readdata,                         --                                         .readdata
			HEX_3_s1_writedata                             => mm_interconnect_0_hex_3_s1_writedata,                        --                                         .writedata
			HEX_3_s1_chipselect                            => mm_interconnect_0_hex_3_s1_chipselect,                       --                                         .chipselect
			HEX_4_s1_address                               => mm_interconnect_0_hex_4_s1_address,                          --                                 HEX_4_s1.address
			HEX_4_s1_write                                 => mm_interconnect_0_hex_4_s1_write,                            --                                         .write
			HEX_4_s1_readdata                              => mm_interconnect_0_hex_4_s1_readdata,                         --                                         .readdata
			HEX_4_s1_writedata                             => mm_interconnect_0_hex_4_s1_writedata,                        --                                         .writedata
			HEX_4_s1_chipselect                            => mm_interconnect_0_hex_4_s1_chipselect,                       --                                         .chipselect
			HEX_5_s1_address                               => mm_interconnect_0_hex_5_s1_address,                          --                                 HEX_5_s1.address
			HEX_5_s1_write                                 => mm_interconnect_0_hex_5_s1_write,                            --                                         .write
			HEX_5_s1_readdata                              => mm_interconnect_0_hex_5_s1_readdata,                         --                                         .readdata
			HEX_5_s1_writedata                             => mm_interconnect_0_hex_5_s1_writedata,                        --                                         .writedata
			HEX_5_s1_chipselect                            => mm_interconnect_0_hex_5_s1_chipselect,                       --                                         .chipselect
			HEX_6_s1_address                               => mm_interconnect_0_hex_6_s1_address,                          --                                 HEX_6_s1.address
			HEX_6_s1_write                                 => mm_interconnect_0_hex_6_s1_write,                            --                                         .write
			HEX_6_s1_readdata                              => mm_interconnect_0_hex_6_s1_readdata,                         --                                         .readdata
			HEX_6_s1_writedata                             => mm_interconnect_0_hex_6_s1_writedata,                        --                                         .writedata
			HEX_6_s1_chipselect                            => mm_interconnect_0_hex_6_s1_chipselect,                       --                                         .chipselect
			HEX_7_s1_address                               => mm_interconnect_0_hex_7_s1_address,                          --                                 HEX_7_s1.address
			HEX_7_s1_write                                 => mm_interconnect_0_hex_7_s1_write,                            --                                         .write
			HEX_7_s1_readdata                              => mm_interconnect_0_hex_7_s1_readdata,                         --                                         .readdata
			HEX_7_s1_writedata                             => mm_interconnect_0_hex_7_s1_writedata,                        --                                         .writedata
			HEX_7_s1_chipselect                            => mm_interconnect_0_hex_7_s1_chipselect,                       --                                         .chipselect
			jtag_uart_0_avalon_jtag_slave_address          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --            jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                         .write
			jtag_uart_0_avalon_jtag_slave_read             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                         .read
			jtag_uart_0_avalon_jtag_slave_readdata         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                         .readdata
			jtag_uart_0_avalon_jtag_slave_writedata        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                         .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                         .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                         .chipselect
			move_left_s1_address                           => mm_interconnect_0_move_left_s1_address,                      --                             move_left_s1.address
			move_left_s1_write                             => mm_interconnect_0_move_left_s1_write,                        --                                         .write
			move_left_s1_readdata                          => mm_interconnect_0_move_left_s1_readdata,                     --                                         .readdata
			move_left_s1_writedata                         => mm_interconnect_0_move_left_s1_writedata,                    --                                         .writedata
			move_left_s1_chipselect                        => mm_interconnect_0_move_left_s1_chipselect,                   --                                         .chipselect
			move_right_s1_address                          => mm_interconnect_0_move_right_s1_address,                     --                            move_right_s1.address
			move_right_s1_write                            => mm_interconnect_0_move_right_s1_write,                       --                                         .write
			move_right_s1_readdata                         => mm_interconnect_0_move_right_s1_readdata,                    --                                         .readdata
			move_right_s1_writedata                        => mm_interconnect_0_move_right_s1_writedata,                   --                                         .writedata
			move_right_s1_chipselect                       => mm_interconnect_0_move_right_s1_chipselect,                  --                                         .chipselect
			nios2_gen2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,      --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,        --                                         .write
			nios2_gen2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,         --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,     --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,    --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,   --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,  --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,  --                                         .debugaccess
			onchip_memory2_0_s1_address                    => mm_interconnect_0_onchip_memory2_0_s1_address,               --                      onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                      => mm_interconnect_0_onchip_memory2_0_s1_write,                 --                                         .write
			onchip_memory2_0_s1_readdata                   => mm_interconnect_0_onchip_memory2_0_s1_readdata,              --                                         .readdata
			onchip_memory2_0_s1_writedata                  => mm_interconnect_0_onchip_memory2_0_s1_writedata,             --                                         .writedata
			onchip_memory2_0_s1_byteenable                 => mm_interconnect_0_onchip_memory2_0_s1_byteenable,            --                                         .byteenable
			onchip_memory2_0_s1_chipselect                 => mm_interconnect_0_onchip_memory2_0_s1_chipselect,            --                                         .chipselect
			onchip_memory2_0_s1_clken                      => mm_interconnect_0_onchip_memory2_0_s1_clken,                 --                                         .clken
			rotate_left_s1_address                         => mm_interconnect_0_rotate_left_s1_address,                    --                           rotate_left_s1.address
			rotate_left_s1_write                           => mm_interconnect_0_rotate_left_s1_write,                      --                                         .write
			rotate_left_s1_readdata                        => mm_interconnect_0_rotate_left_s1_readdata,                   --                                         .readdata
			rotate_left_s1_writedata                       => mm_interconnect_0_rotate_left_s1_writedata,                  --                                         .writedata
			rotate_left_s1_chipselect                      => mm_interconnect_0_rotate_left_s1_chipselect,                 --                                         .chipselect
			rotate_right_s1_address                        => mm_interconnect_0_rotate_right_s1_address,                   --                          rotate_right_s1.address
			rotate_right_s1_write                          => mm_interconnect_0_rotate_right_s1_write,                     --                                         .write
			rotate_right_s1_readdata                       => mm_interconnect_0_rotate_right_s1_readdata,                  --                                         .readdata
			rotate_right_s1_writedata                      => mm_interconnect_0_rotate_right_s1_writedata,                 --                                         .writedata
			rotate_right_s1_chipselect                     => mm_interconnect_0_rotate_right_s1_chipselect,                --                                         .chipselect
			row_0_s1_address                               => mm_interconnect_0_row_0_s1_address,                          --                                 row_0_s1.address
			row_0_s1_write                                 => mm_interconnect_0_row_0_s1_write,                            --                                         .write
			row_0_s1_readdata                              => mm_interconnect_0_row_0_s1_readdata,                         --                                         .readdata
			row_0_s1_writedata                             => mm_interconnect_0_row_0_s1_writedata,                        --                                         .writedata
			row_0_s1_chipselect                            => mm_interconnect_0_row_0_s1_chipselect,                       --                                         .chipselect
			row_1_s1_address                               => mm_interconnect_0_row_1_s1_address,                          --                                 row_1_s1.address
			row_1_s1_write                                 => mm_interconnect_0_row_1_s1_write,                            --                                         .write
			row_1_s1_readdata                              => mm_interconnect_0_row_1_s1_readdata,                         --                                         .readdata
			row_1_s1_writedata                             => mm_interconnect_0_row_1_s1_writedata,                        --                                         .writedata
			row_1_s1_chipselect                            => mm_interconnect_0_row_1_s1_chipselect,                       --                                         .chipselect
			row_10_s1_address                              => mm_interconnect_0_row_10_s1_address,                         --                                row_10_s1.address
			row_10_s1_write                                => mm_interconnect_0_row_10_s1_write,                           --                                         .write
			row_10_s1_readdata                             => mm_interconnect_0_row_10_s1_readdata,                        --                                         .readdata
			row_10_s1_writedata                            => mm_interconnect_0_row_10_s1_writedata,                       --                                         .writedata
			row_10_s1_chipselect                           => mm_interconnect_0_row_10_s1_chipselect,                      --                                         .chipselect
			row_11_s1_address                              => mm_interconnect_0_row_11_s1_address,                         --                                row_11_s1.address
			row_11_s1_write                                => mm_interconnect_0_row_11_s1_write,                           --                                         .write
			row_11_s1_readdata                             => mm_interconnect_0_row_11_s1_readdata,                        --                                         .readdata
			row_11_s1_writedata                            => mm_interconnect_0_row_11_s1_writedata,                       --                                         .writedata
			row_11_s1_chipselect                           => mm_interconnect_0_row_11_s1_chipselect,                      --                                         .chipselect
			row_12_s1_address                              => mm_interconnect_0_row_12_s1_address,                         --                                row_12_s1.address
			row_12_s1_write                                => mm_interconnect_0_row_12_s1_write,                           --                                         .write
			row_12_s1_readdata                             => mm_interconnect_0_row_12_s1_readdata,                        --                                         .readdata
			row_12_s1_writedata                            => mm_interconnect_0_row_12_s1_writedata,                       --                                         .writedata
			row_12_s1_chipselect                           => mm_interconnect_0_row_12_s1_chipselect,                      --                                         .chipselect
			row_13_s1_address                              => mm_interconnect_0_row_13_s1_address,                         --                                row_13_s1.address
			row_13_s1_write                                => mm_interconnect_0_row_13_s1_write,                           --                                         .write
			row_13_s1_readdata                             => mm_interconnect_0_row_13_s1_readdata,                        --                                         .readdata
			row_13_s1_writedata                            => mm_interconnect_0_row_13_s1_writedata,                       --                                         .writedata
			row_13_s1_chipselect                           => mm_interconnect_0_row_13_s1_chipselect,                      --                                         .chipselect
			row_14_s1_address                              => mm_interconnect_0_row_14_s1_address,                         --                                row_14_s1.address
			row_14_s1_write                                => mm_interconnect_0_row_14_s1_write,                           --                                         .write
			row_14_s1_readdata                             => mm_interconnect_0_row_14_s1_readdata,                        --                                         .readdata
			row_14_s1_writedata                            => mm_interconnect_0_row_14_s1_writedata,                       --                                         .writedata
			row_14_s1_chipselect                           => mm_interconnect_0_row_14_s1_chipselect,                      --                                         .chipselect
			row_15_s1_address                              => mm_interconnect_0_row_15_s1_address,                         --                                row_15_s1.address
			row_15_s1_write                                => mm_interconnect_0_row_15_s1_write,                           --                                         .write
			row_15_s1_readdata                             => mm_interconnect_0_row_15_s1_readdata,                        --                                         .readdata
			row_15_s1_writedata                            => mm_interconnect_0_row_15_s1_writedata,                       --                                         .writedata
			row_15_s1_chipselect                           => mm_interconnect_0_row_15_s1_chipselect,                      --                                         .chipselect
			row_16_s1_address                              => mm_interconnect_0_row_16_s1_address,                         --                                row_16_s1.address
			row_16_s1_write                                => mm_interconnect_0_row_16_s1_write,                           --                                         .write
			row_16_s1_readdata                             => mm_interconnect_0_row_16_s1_readdata,                        --                                         .readdata
			row_16_s1_writedata                            => mm_interconnect_0_row_16_s1_writedata,                       --                                         .writedata
			row_16_s1_chipselect                           => mm_interconnect_0_row_16_s1_chipselect,                      --                                         .chipselect
			row_17_s1_address                              => mm_interconnect_0_row_17_s1_address,                         --                                row_17_s1.address
			row_17_s1_write                                => mm_interconnect_0_row_17_s1_write,                           --                                         .write
			row_17_s1_readdata                             => mm_interconnect_0_row_17_s1_readdata,                        --                                         .readdata
			row_17_s1_writedata                            => mm_interconnect_0_row_17_s1_writedata,                       --                                         .writedata
			row_17_s1_chipselect                           => mm_interconnect_0_row_17_s1_chipselect,                      --                                         .chipselect
			row_18_s1_address                              => mm_interconnect_0_row_18_s1_address,                         --                                row_18_s1.address
			row_18_s1_write                                => mm_interconnect_0_row_18_s1_write,                           --                                         .write
			row_18_s1_readdata                             => mm_interconnect_0_row_18_s1_readdata,                        --                                         .readdata
			row_18_s1_writedata                            => mm_interconnect_0_row_18_s1_writedata,                       --                                         .writedata
			row_18_s1_chipselect                           => mm_interconnect_0_row_18_s1_chipselect,                      --                                         .chipselect
			row_19_s1_address                              => mm_interconnect_0_row_19_s1_address,                         --                                row_19_s1.address
			row_19_s1_write                                => mm_interconnect_0_row_19_s1_write,                           --                                         .write
			row_19_s1_readdata                             => mm_interconnect_0_row_19_s1_readdata,                        --                                         .readdata
			row_19_s1_writedata                            => mm_interconnect_0_row_19_s1_writedata,                       --                                         .writedata
			row_19_s1_chipselect                           => mm_interconnect_0_row_19_s1_chipselect,                      --                                         .chipselect
			row_2_s1_address                               => mm_interconnect_0_row_2_s1_address,                          --                                 row_2_s1.address
			row_2_s1_write                                 => mm_interconnect_0_row_2_s1_write,                            --                                         .write
			row_2_s1_readdata                              => mm_interconnect_0_row_2_s1_readdata,                         --                                         .readdata
			row_2_s1_writedata                             => mm_interconnect_0_row_2_s1_writedata,                        --                                         .writedata
			row_2_s1_chipselect                            => mm_interconnect_0_row_2_s1_chipselect,                       --                                         .chipselect
			row_20_s1_address                              => mm_interconnect_0_row_20_s1_address,                         --                                row_20_s1.address
			row_20_s1_write                                => mm_interconnect_0_row_20_s1_write,                           --                                         .write
			row_20_s1_readdata                             => mm_interconnect_0_row_20_s1_readdata,                        --                                         .readdata
			row_20_s1_writedata                            => mm_interconnect_0_row_20_s1_writedata,                       --                                         .writedata
			row_20_s1_chipselect                           => mm_interconnect_0_row_20_s1_chipselect,                      --                                         .chipselect
			row_21_s1_address                              => mm_interconnect_0_row_21_s1_address,                         --                                row_21_s1.address
			row_21_s1_write                                => mm_interconnect_0_row_21_s1_write,                           --                                         .write
			row_21_s1_readdata                             => mm_interconnect_0_row_21_s1_readdata,                        --                                         .readdata
			row_21_s1_writedata                            => mm_interconnect_0_row_21_s1_writedata,                       --                                         .writedata
			row_21_s1_chipselect                           => mm_interconnect_0_row_21_s1_chipselect,                      --                                         .chipselect
			row_22_s1_address                              => mm_interconnect_0_row_22_s1_address,                         --                                row_22_s1.address
			row_22_s1_write                                => mm_interconnect_0_row_22_s1_write,                           --                                         .write
			row_22_s1_readdata                             => mm_interconnect_0_row_22_s1_readdata,                        --                                         .readdata
			row_22_s1_writedata                            => mm_interconnect_0_row_22_s1_writedata,                       --                                         .writedata
			row_22_s1_chipselect                           => mm_interconnect_0_row_22_s1_chipselect,                      --                                         .chipselect
			row_23_s1_address                              => mm_interconnect_0_row_23_s1_address,                         --                                row_23_s1.address
			row_23_s1_write                                => mm_interconnect_0_row_23_s1_write,                           --                                         .write
			row_23_s1_readdata                             => mm_interconnect_0_row_23_s1_readdata,                        --                                         .readdata
			row_23_s1_writedata                            => mm_interconnect_0_row_23_s1_writedata,                       --                                         .writedata
			row_23_s1_chipselect                           => mm_interconnect_0_row_23_s1_chipselect,                      --                                         .chipselect
			row_3_s1_address                               => mm_interconnect_0_row_3_s1_address,                          --                                 row_3_s1.address
			row_3_s1_write                                 => mm_interconnect_0_row_3_s1_write,                            --                                         .write
			row_3_s1_readdata                              => mm_interconnect_0_row_3_s1_readdata,                         --                                         .readdata
			row_3_s1_writedata                             => mm_interconnect_0_row_3_s1_writedata,                        --                                         .writedata
			row_3_s1_chipselect                            => mm_interconnect_0_row_3_s1_chipselect,                       --                                         .chipselect
			row_4_s1_address                               => mm_interconnect_0_row_4_s1_address,                          --                                 row_4_s1.address
			row_4_s1_write                                 => mm_interconnect_0_row_4_s1_write,                            --                                         .write
			row_4_s1_readdata                              => mm_interconnect_0_row_4_s1_readdata,                         --                                         .readdata
			row_4_s1_writedata                             => mm_interconnect_0_row_4_s1_writedata,                        --                                         .writedata
			row_4_s1_chipselect                            => mm_interconnect_0_row_4_s1_chipselect,                       --                                         .chipselect
			row_5_s1_address                               => mm_interconnect_0_row_5_s1_address,                          --                                 row_5_s1.address
			row_5_s1_write                                 => mm_interconnect_0_row_5_s1_write,                            --                                         .write
			row_5_s1_readdata                              => mm_interconnect_0_row_5_s1_readdata,                         --                                         .readdata
			row_5_s1_writedata                             => mm_interconnect_0_row_5_s1_writedata,                        --                                         .writedata
			row_5_s1_chipselect                            => mm_interconnect_0_row_5_s1_chipselect,                       --                                         .chipselect
			row_6_s1_address                               => mm_interconnect_0_row_6_s1_address,                          --                                 row_6_s1.address
			row_6_s1_write                                 => mm_interconnect_0_row_6_s1_write,                            --                                         .write
			row_6_s1_readdata                              => mm_interconnect_0_row_6_s1_readdata,                         --                                         .readdata
			row_6_s1_writedata                             => mm_interconnect_0_row_6_s1_writedata,                        --                                         .writedata
			row_6_s1_chipselect                            => mm_interconnect_0_row_6_s1_chipselect,                       --                                         .chipselect
			row_7_s1_address                               => mm_interconnect_0_row_7_s1_address,                          --                                 row_7_s1.address
			row_7_s1_write                                 => mm_interconnect_0_row_7_s1_write,                            --                                         .write
			row_7_s1_readdata                              => mm_interconnect_0_row_7_s1_readdata,                         --                                         .readdata
			row_7_s1_writedata                             => mm_interconnect_0_row_7_s1_writedata,                        --                                         .writedata
			row_7_s1_chipselect                            => mm_interconnect_0_row_7_s1_chipselect,                       --                                         .chipselect
			row_8_s1_address                               => mm_interconnect_0_row_8_s1_address,                          --                                 row_8_s1.address
			row_8_s1_write                                 => mm_interconnect_0_row_8_s1_write,                            --                                         .write
			row_8_s1_readdata                              => mm_interconnect_0_row_8_s1_readdata,                         --                                         .readdata
			row_8_s1_writedata                             => mm_interconnect_0_row_8_s1_writedata,                        --                                         .writedata
			row_8_s1_chipselect                            => mm_interconnect_0_row_8_s1_chipselect,                       --                                         .chipselect
			row_9_s1_address                               => mm_interconnect_0_row_9_s1_address,                          --                                 row_9_s1.address
			row_9_s1_write                                 => mm_interconnect_0_row_9_s1_write,                            --                                         .write
			row_9_s1_readdata                              => mm_interconnect_0_row_9_s1_readdata,                         --                                         .readdata
			row_9_s1_writedata                             => mm_interconnect_0_row_9_s1_writedata,                        --                                         .writedata
			row_9_s1_chipselect                            => mm_interconnect_0_row_9_s1_chipselect,                       --                                         .chipselect
			sram_0_avalon_sram_slave_address               => mm_interconnect_0_sram_0_avalon_sram_slave_address,          --                 sram_0_avalon_sram_slave.address
			sram_0_avalon_sram_slave_write                 => mm_interconnect_0_sram_0_avalon_sram_slave_write,            --                                         .write
			sram_0_avalon_sram_slave_read                  => mm_interconnect_0_sram_0_avalon_sram_slave_read,             --                                         .read
			sram_0_avalon_sram_slave_readdata              => mm_interconnect_0_sram_0_avalon_sram_slave_readdata,         --                                         .readdata
			sram_0_avalon_sram_slave_writedata             => mm_interconnect_0_sram_0_avalon_sram_slave_writedata,        --                                         .writedata
			sram_0_avalon_sram_slave_byteenable            => mm_interconnect_0_sram_0_avalon_sram_slave_byteenable,       --                                         .byteenable
			sram_0_avalon_sram_slave_readdatavalid         => mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid     --                                         .readdatavalid
		);

	irq_mapper : component sram_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,       -- receiver5.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_row_0_s1_write_ports_inv <= not mm_interconnect_0_row_0_s1_write;

	mm_interconnect_0_row_1_s1_write_ports_inv <= not mm_interconnect_0_row_1_s1_write;

	mm_interconnect_0_row_2_s1_write_ports_inv <= not mm_interconnect_0_row_2_s1_write;

	mm_interconnect_0_row_3_s1_write_ports_inv <= not mm_interconnect_0_row_3_s1_write;

	mm_interconnect_0_row_4_s1_write_ports_inv <= not mm_interconnect_0_row_4_s1_write;

	mm_interconnect_0_row_5_s1_write_ports_inv <= not mm_interconnect_0_row_5_s1_write;

	mm_interconnect_0_row_6_s1_write_ports_inv <= not mm_interconnect_0_row_6_s1_write;

	mm_interconnect_0_row_7_s1_write_ports_inv <= not mm_interconnect_0_row_7_s1_write;

	mm_interconnect_0_row_8_s1_write_ports_inv <= not mm_interconnect_0_row_8_s1_write;

	mm_interconnect_0_row_9_s1_write_ports_inv <= not mm_interconnect_0_row_9_s1_write;

	mm_interconnect_0_row_11_s1_write_ports_inv <= not mm_interconnect_0_row_11_s1_write;

	mm_interconnect_0_row_12_s1_write_ports_inv <= not mm_interconnect_0_row_12_s1_write;

	mm_interconnect_0_row_13_s1_write_ports_inv <= not mm_interconnect_0_row_13_s1_write;

	mm_interconnect_0_row_14_s1_write_ports_inv <= not mm_interconnect_0_row_14_s1_write;

	mm_interconnect_0_row_15_s1_write_ports_inv <= not mm_interconnect_0_row_15_s1_write;

	mm_interconnect_0_row_16_s1_write_ports_inv <= not mm_interconnect_0_row_16_s1_write;

	mm_interconnect_0_row_17_s1_write_ports_inv <= not mm_interconnect_0_row_17_s1_write;

	mm_interconnect_0_row_18_s1_write_ports_inv <= not mm_interconnect_0_row_18_s1_write;

	mm_interconnect_0_row_19_s1_write_ports_inv <= not mm_interconnect_0_row_19_s1_write;

	mm_interconnect_0_row_20_s1_write_ports_inv <= not mm_interconnect_0_row_20_s1_write;

	mm_interconnect_0_row_21_s1_write_ports_inv <= not mm_interconnect_0_row_21_s1_write;

	mm_interconnect_0_row_22_s1_write_ports_inv <= not mm_interconnect_0_row_22_s1_write;

	mm_interconnect_0_row_23_s1_write_ports_inv <= not mm_interconnect_0_row_23_s1_write;

	mm_interconnect_0_row_10_s1_write_ports_inv <= not mm_interconnect_0_row_10_s1_write;

	mm_interconnect_0_move_left_s1_write_ports_inv <= not mm_interconnect_0_move_left_s1_write;

	mm_interconnect_0_move_right_s1_write_ports_inv <= not mm_interconnect_0_move_right_s1_write;

	mm_interconnect_0_rotate_left_s1_write_ports_inv <= not mm_interconnect_0_rotate_left_s1_write;

	mm_interconnect_0_rotate_right_s1_write_ports_inv <= not mm_interconnect_0_rotate_right_s1_write;

	mm_interconnect_0_frame_timer_s1_write_ports_inv <= not mm_interconnect_0_frame_timer_s1_write;

	mm_interconnect_0_hex_0_s1_write_ports_inv <= not mm_interconnect_0_hex_0_s1_write;

	mm_interconnect_0_hex_1_s1_write_ports_inv <= not mm_interconnect_0_hex_1_s1_write;

	mm_interconnect_0_hex_2_s1_write_ports_inv <= not mm_interconnect_0_hex_2_s1_write;

	mm_interconnect_0_hex_3_s1_write_ports_inv <= not mm_interconnect_0_hex_3_s1_write;

	mm_interconnect_0_hex_4_s1_write_ports_inv <= not mm_interconnect_0_hex_4_s1_write;

	mm_interconnect_0_hex_5_s1_write_ports_inv <= not mm_interconnect_0_hex_5_s1_write;

	mm_interconnect_0_hex_6_s1_write_ports_inv <= not mm_interconnect_0_hex_6_s1_write;

	mm_interconnect_0_hex_7_s1_write_ports_inv <= not mm_interconnect_0_hex_7_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of sram
